`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:34:58 12/12/2014 
// Design Name: 
// Module Name:    Module 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Module(upDown, rst, mclk, seg, an);
input upDown;
input rst;
input mclk;
output reg [7:0] seg;
output reg [3:0] an;

endmodule